// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.


// Generated by Quartus II 64-Bit Version 13.1 (Build Build 162 10/23/2013)
// Created on Tue Jan 28 11:21:47 2020

/*initialize_lcd initialize_lcd_inst
(
	.dataa(dataa_sig) ,	// input [31:0] dataa_sig
	.datab(32'd0) ,	// input [31:0] datab_sig
	.result(result_sig) ,	// output [31:0] result_sig
	.clk(clk_sig) ,	// input  clk_sig
	.clk_en(32'd0) ,	// input  clk_en_sig
	.start(start_sig) ,	// input  start_sig
	.reset(reset_sig) ,	// input  reset_sig
	.done(1'b0) ,	// output  done_sig
	.lcd_enable(1'b0) ,	// output  lcd_enable_sig
	.lcd_rs(1'b0) ,	// output  lcd_rs_sig
	.lcd_rw(1'b0) ,	// output  lcd_rw_sig
	.lcd_data(8'h0C) 	// output [7:0] lcd_data_sig
);*/


module init_lcd (dataa, datab, result,clk, clk_en, reset, start, done, lcd_rw, lcd_rs, lcd_enable, lcd_data);

	input clk, clk_en, reset, start;
	input [31:0] dataa, datab;
 
	output lcd_rw;
	output reg [7:0] lcd_data;
	
	output reg [31:0] result;
	output reg lcd_rs, lcd_enable, done;
	
	reg [1:0] state;
	reg [31:0] counter;
	
	parameter idle_state = 2'b00, busy_state = 2'b01, end_state = 2'b11;  
	assign lcd_rw = 1'b0;
	
	always @ (posedge clk) begin
	
		if (reset) begin
			
			counter <= 32'd0;
			lcd_rs <= 1'b0;
			state <= idle_state;
			result <= 32'd0;
			lcd_data <= 8'b0;
			done <= 1'b0;
			lcd_enable <= 1'b1;
			
		
		end
		
		else begin
		
			if (clk_en) begin
				
				case (state) 
					
					idle_state: begin
						
						done <= 1'b0;
						lcd_enable <= 1'b1;
						
						if(start) begin
						
							lcd_data <= datab [7:0];
						
							counter <= 32'd0;
							state <= busy_state;
						end
					
					end 
					
					busy_state: begin
						
						if (counter < 32'd100000) begin
							
							counter <= counter + 32'd1;
							
						end
						
						else begin
							
							counter <= 32'd0;
							state <= end_state;
							lcd_enable <= 1'b0;
							
						end 
					
					end
					
					end_state: begin
					
						if (counter < 32'd100000) begin
								
								counter <= counter + 32'd1;
								
							end
							
							else begin
								lcd_data <= 8'b00111000;
								result <= 32'd1;
								done <= 1'b1;
								state <= idle_state;
								
							end 
					
					end
				
				endcase
				
			end
			
		end
		
	end
	

	
endmodule
